VERSION 5.8 ;

BUSBITCHARS "[]" ;

DIVIDERCHAR "/" ;

UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.000500 ;

CLEARANCEMEASURE EUCLIDEAN ;
USEMINSPACING OBS ON ;

SITE CoreSite
    CLASS CORE ;
    SIZE 0.200000 BY 1.710000 ; 
END CoreSite

LAYER Metal1
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    MINWIDTH 0.060000 ;
    AREA 0.020000 ;
    WIDTH 0.060000 ;
    SPACING 0.060000 ;
    SPACING 0.090000 ENDOFLINE 0.090000 WITHIN 0.025000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.060000
      WIDTH  0.100000  0.100000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 0.190000 0.190000 ;
END Metal1

LAYER Via1
    TYPE CUT ;
    SPACING 0.070000 ;
    WIDTH 0.06 ;
END Via1

LAYER Metal2
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    MINWIDTH 0.070000 ;
    AREA 0.020000 ;
    WIDTH 0.070000 ;
    SPACING 0.070000 ;
    SPACING 0.100000 ENDOFLINE 0.100000 WITHIN 0.035000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.070000
      WIDTH  0.100000  0.150000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 0.200000 0.200000 ;
END Metal2

LAYER Via2
    TYPE CUT ;
    SPACING 0.070000 ;
    WIDTH 0.07 ;
END Via2

LAYER Metal3
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    MINWIDTH 0.070000 ;
    AREA 0.020000 ;
    WIDTH 0.070000 ;
    SPACING 0.070000 ;
    SPACING 0.100000 ENDOFLINE 0.100000 WITHIN 0.035000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.070000
      WIDTH  0.100000  0.150000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 0.200000 0.200000 ;
END Metal3

LAYER Via3
    TYPE CUT ;
    SPACING 0.070000 ;
    WIDTH 0.07 ;
END Via3

LAYER Metal4
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    MINWIDTH 0.070000 ;
    AREA 0.020000 ;
    WIDTH 0.070000 ;
    SPACING 0.070000 ;
    SPACING 0.100000 ENDOFLINE 0.100000 WITHIN 0.035000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.070000
      WIDTH  0.100000  0.150000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 0.200000 0.200000 ;
END Metal4

LAYER Via4
    TYPE CUT ;
    SPACING 0.070000 ;
    WIDTH 0.07 ;
END Via4

LAYER Metal5
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    MINWIDTH 0.070000 ;
    AREA 0.020000 ;
    WIDTH 0.070000 ;
    SPACING 0.070000 ;
    SPACING 0.100000 ENDOFLINE 0.100000 WITHIN 0.035000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.070000
      WIDTH  0.100000  0.150000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 0.200000 0.200000 ;
END Metal5

LAYER Via5
    TYPE CUT ;
    SPACING 0.070000 ;
    WIDTH 0.07 ;
END Via5

LAYER Metal6
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    MINWIDTH 0.070000 ;
    AREA 0.020000 ;
    WIDTH 0.070000 ;
    SPACING 0.070000 ;
    SPACING 0.100000 ENDOFLINE 0.100000 WITHIN 0.035000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.070000
      WIDTH  0.100000  0.150000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 0.200000 0.200000 ;
END Metal6

LAYER Via6
    TYPE CUT ;
    SPACING 0.070000 ;
    WIDTH 0.07 ;
END Via6

LAYER Metal7
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    MINWIDTH 0.070000 ;
    AREA 0.020000 ;
    WIDTH 0.070000 ;
    SPACING 0.070000 ;
    SPACING 0.100000 ENDOFLINE 0.100000 WITHIN 0.035000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.070000
      WIDTH  0.100000  0.150000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 0.200000 0.200000 ;
END Metal7

LAYER Via7
    TYPE CUT ;
    SPACING 0.070000 ;
    WIDTH 0.07 ;
END Via7

LAYER Metal8
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    MINWIDTH 0.070000 ;
    AREA 0.020000 ;
    WIDTH 0.070000 ;
    SPACING 0.070000 ;
    SPACING 0.100000 ENDOFLINE 0.100000 WITHIN 0.035000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.070000
      WIDTH  0.100000  0.150000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 0.200000 0.200000 ;
END Metal8

LAYER Via8
    TYPE CUT ;
    SPACING 0.070000 ;
    WIDTH 0.07 ;
END Via8

LAYER Metal9
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    MINWIDTH 0.070000 ;
    AREA 0.020000 ;
    WIDTH 0.070000 ;
    SPACING 0.070000 ;
    SPACING 0.100000 ENDOFLINE 0.100000 WITHIN 0.035000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.070000
      WIDTH  0.100000  0.150000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 0.330000 0.330000 ;
END Metal9

LAYER OVERLAP
    TYPE OVERLAP ;
END OVERLAP

VIA VIA12_1C DEFAULT 
    LAYER Metal1 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via1 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal2 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA12_1C

VIA VIA12_1C_H DEFAULT 
    LAYER Metal1 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via1 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal2 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA12_1C_H

VIA VIA12_1C_V DEFAULT 
    LAYER Metal1 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via1 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal2 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA12_1C_V

VIA VIA23_1C DEFAULT 
    LAYER Metal2 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA23_1C

VIA VIA23_1C_H DEFAULT 
    LAYER Metal2 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA23_1C_H

VIA VIA23_1C_V DEFAULT 
    LAYER Metal2 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal3 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA23_1C_V

VIA VIA23_1ST_N DEFAULT 
    LAYER Metal2 ;
        RECT -0.035000 -0.065000 0.035000 0.325000 ;
    LAYER Via2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA23_1ST_N

VIA VIA23_1ST_S DEFAULT 
    LAYER Metal2 ;
        RECT -0.035000 -0.325000 0.035000 0.065000 ;
    LAYER Via2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA23_1ST_S

VIA VIA34_1C DEFAULT 
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA34_1C

VIA VIA34_1C_H DEFAULT 
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal4 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA34_1C_H

VIA VIA34_1C_V DEFAULT 
    LAYER Metal3 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA34_1C_V

VIA VIA34_1ST_E DEFAULT 
    LAYER Metal3 ;
        RECT -0.065000 -0.035000 0.325000 0.035000 ;
    LAYER Via3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA34_1ST_E

VIA VIA34_1ST_W DEFAULT 
    LAYER Metal3 ;
        RECT -0.325000 -0.035000 0.065000 0.035000 ;
    LAYER Via3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA34_1ST_W

VIA VIA45_1C DEFAULT 
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal5 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA45_1C

VIA VIA45_1C_H DEFAULT 
    LAYER Metal4 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal5 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA45_1C_H

VIA VIA45_1C_V DEFAULT 
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal5 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA45_1C_V

VIA VIA45_1ST_N DEFAULT 
    LAYER Metal4 ;
        RECT -0.035000 -0.065000 0.035000 0.325000 ;
    LAYER Via4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal5 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA45_1ST_N

VIA VIA45_1ST_S DEFAULT 
    LAYER Metal4 ;
        RECT -0.035000 -0.325000 0.035000 0.065000 ;
    LAYER Via4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal5 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA45_1ST_S

VIA VIA5_0_VH DEFAULT 
    LAYER Metal5 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via5 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal6 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA5_0_VH

VIA VIA6_0_HV DEFAULT 
    LAYER Metal6 ;
        RECT -0.260000 -0.200000 0.260000 0.200000 ;
    LAYER Via6 ;
        RECT -0.180000 -0.180000 0.180000 0.180000 ;
    LAYER Metal7 ;
        RECT -0.200000 -0.260000 0.200000 0.260000 ;
END VIA6_0_HV

VIA VIA7_0_VH DEFAULT 
    LAYER Metal7 ;
        RECT -0.200000 -0.260000 0.200000 0.260000 ;
    LAYER Via7 ;
        RECT -0.180000 -0.180000 0.180000 0.180000 ;
    LAYER Metal8 ;
        RECT -0.260000 -0.200000 0.260000 0.200000 ;
END VIA7_0_VH

VIA VIA8_0_VH DEFAULT 
    LAYER Metal8 ;
        RECT -0.200000 -0.260000 0.200000 0.260000 ;
    LAYER Via8 ;
        RECT -0.180000 -0.180000 0.180000 0.180000 ;
    LAYER Metal9 ;
        RECT -0.260000 -0.200000 0.260000 0.200000 ;
END VIA8_0_VH


MACRO AOI221X2
    CLASS CORE ;
    FOREIGN AOI221X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.600000 BY 1.710000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.235000 0.625000 0.365000 0.715000 ;
        RECT 0.285000 0.610000 0.960000 0.690000 ;
        RECT 0.285000 0.610000 0.365000 0.715000 ;
        RECT 0.235000 0.625000 0.960000 0.690000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.660000 0.765000 0.740000 1.065000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.635000 0.625000 1.765000 0.715000 ;
        RECT 1.240000 0.635000 1.935000 0.715000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.435000 0.815000 1.935000 0.895000 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.065000 0.815000 2.565000 0.895000 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.650000 2.600000 1.710000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 0.000000 2.600000 0.060000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.060000 0.790000 1.140000 0.920000 ;
        RECT 2.220000 0.995000 2.280000 1.135000 ;
        RECT 1.080000 0.995000 2.280000 1.055000 ;
        RECT 1.080000 0.450000 1.140000 1.055000 ;
        RECT 0.605000 0.450000 2.170000 0.510000 ;
        END
    END Y
END AOI221X2

MACRO NAND3X2
    CLASS CORE ;
    FOREIGN NAND3X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.600000 BY 1.710000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.260000 0.600000 0.370000 0.735000 ;
        RECT 1.240000 0.495000 1.300000 0.735000 ;
        RECT 0.310000 0.495000 1.300000 0.555000 ;
        RECT 0.310000 0.495000 0.370000 0.735000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.060000 0.655000 1.140000 0.920000 ;
        RECT 0.470000 0.655000 1.140000 0.715000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.520000 0.815000 0.765000 0.955000 ;
        RECT 0.520000 0.815000 0.960000 0.895000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.650000 1.600000 1.710000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 0.000000 1.600000 0.060000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.435000 1.005000 1.565000 1.115000 ;
        RECT 0.360000 1.055000 0.430000 1.335000 ;
        RECT 1.505000 0.335000 1.565000 1.115000 ;
        RECT 1.190000 1.055000 1.250000 1.335000 ;
        RECT 0.795000 0.335000 1.565000 0.395000 ;
        RECT 0.780000 1.055000 0.840000 1.335000 ;
        RECT 0.360000 1.055000 1.565000 1.115000 ;
        END
    END Y
END NAND3X2

END LIBRARY
